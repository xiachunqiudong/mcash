// CROSS BAR
bind spw_buffer spw_buffer_assert #(.PTR_WIDTH(3)) u_spw_buffer_assert (.*);
bind cross_bar_top cross_bar_assert u_cross_bar_assert(.*);
bind cross_bar_rob cross_bar_rob_assert u_cross_bar_rob_assert(.*);