`define WBUFFER_AW
`define FREELIST_WIDTH 1 << WBUFFER_AW